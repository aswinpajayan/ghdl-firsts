library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.Numeric_Std.all;

entity Imem is
    Port ( address : in  STD_LOGIC_VECTOR (15 downto 0);
           data_out : out  STD_LOGIC_VECTOR (15 downto 0));
end Imem;

architecture arc_Imem of Imem is

type memory16 is array (0 to (2**16)-1) of STD_LOGIC_VECTOR (15 downto 0);

signal memory : memory16 := 
(
--  X"FFFF",	
   B"0000_001_010_111_000", --R7 = 0
--    X"0000",
	X"FFFF",	
	B"0110_110_0_00011111",	--LM R1
	B"0000_001_010_011_000", -- ADD R3,R1,R2 ---- 12=3+9
	B"0010_011_100_000_000", -- NDU R0,R3,R4 ---- R0 =0000 0000 0000 1100 nand 0000 0000 0001 1010 = 1111 1111 1111 0111 
	B"0000_011_000_001_001", -- ADZ R1,R3,R0 ---- R1 = 9 (Write signal zero) but carry flag was modified
	B"0000_001_011_101_010", -- ADC R5,R1,R3 ---- 21 = 9+12
	B"0000_001_011_101_010", -- ADC R5,R1,R3 ---- 21 = 9+12 Cy for last zero (Write signal zero)
	B"1000_110_000000000",  --JAL R6,0 --halt


    B"0110_110_0_00011111",	--LM R1
--    B"0101_000_110_000000",	--SW R0,R6,0
--    B"0110_110_0_00100000",	--LM R6
--    B"0000_000_001_010_000", -- ADD R2,R0,R1 ----17=8+9
    B"0000_001_010_011_000", -- ADD R3,R1,R2 ---- 12=3+9
    B"0010_011_100_000_000", -- NDU R0,R3,R4 ---- R0 =0000 0000 0000 1100 nand 0000 0000 0001 1010 = 1111 1111 1111 0111 
    B"0000_011_000_001_001", -- ADZ R1,R3,R0 ---- R1 = 9 but carry flag was modified
    B"0000_001_011_101_010", -- ADC R5,R1,R3 ---- 21 = 9+12
    B"0000_001_011_101_010", -- ADC R5,R1,R3 ---- 21 = 9+12
--    B"1100_011_100_000010",	--BEQ R3,R4,000002
--    B"0000_011_010_100_000", -- ADD R4,R3,R2 ----43=26+17  
--    B"0000_011_010_100_000", -- ADD R4,R3,R2 ----43=26+17 
--    B"0000_011_010_100_000", -- ADD R4,R3,R2 ----43=26+17 
--    B"0110_110_0_10000001",	--LM R6          
--    B"0100_100_110_000001", --LW R4,R6,1;
--    B"0100_101_110_000001", --LW R4,R6,0;
--    B"0000_010_011_000_000", -- ADD R0,R3,R2 ----43=26+17
--    B"0000_010_011_000_000", -- ADD R0,R3,R2 ----43=26+17
--    B"0000_100_010_101_000", -- ADD R5,R4,R2 ----60=43+17 43=26+17 26=9+17
--    B"0100_111_110_000001", --LW R7,R6,1;
--    B"0011_111_000000000", --LHI R7,3; 
--    B"0100_100_110_000000", --LW R4,R6,0;               
--    B"0100_101_110_000001", --LW R5,R6,1;
--    B"0000_101_110_111_000", -- ADD R7,R6,R1 ----9=0+9
--    B"0000_000_001_010_010", -- ADC R2,R0,R1 ----17=8+9     --8+65534=6
--    B"0000_001_010_011_010", -- ADC R3,R1,R2 ----12=9+3     --65534+3=1
--    B"0000_011_010_100_010", -- ADC R4,R3,R2 ----11=8+3     --1+3=4
--    B"0000_100_011_101_010", -- ADC R5,R4,R3 ----8=0+8      --4+1=5
--    B"0010_000_001_010_001", -- NDZ R2,R0,R1 
--    B"0010_001_010_011_001", -- NDZ R3,R1,R2 
--    B"0010_011_010_100_001", -- NDZ R4,R3,R2 
--    B"0010_100_011_101_001", -- NDZ R5,R4,R3 
--    B"0001_000_010_000010", -- ADI R2,R0,000010 --8+2=10
--    B"0001_001_011_000100", -- ADI R3,R1,000100 --65534+4=2
--    B"1001_100_001_000000",	--JLR R4,R1
--    B"0001_011_100_001010", -- ADI R4,R3,001010 --2+10=12
--    B"0001_100_101_110011", -- ADI R5,R4,110011 --12+  
--    B"0101_000_110_000000",	--SW R0,R6,0
--    B"0101_000_110_000000",	--SW R0,R6,0
    B"1000_110_000000000",  --JAL R6,0 --halt   
--    B"0000_000_001_010_000", -- ADD R2,R0,R1
--    B"0000_001_010_011_000", -- ADD R3,R1,R2 
--    B"1000_110_000000000",  --JAL R6,0 --halt
--    B"0011_000_000000001", --LHI R1,1;
--    B"0011_001_000000010", --LHI R2,2;
--    B"0011_010_000000011", --LHI R3,3;
    B"0011_111_000000011", --LHI R7,3; 
	B"1001_101_100_000000",	--JLR
	B"0001_010_001_000000",	--ADI
	B"1001_101_100_000000",	--JLR
	B"0001_011_001_000000",	--ADI
	B"1001_101_100_000000",	--JLR
	B"0010_000_001_000_000",--NDU
	B"1100_100_101_000010",	--BEQ
	B"0001_101_111_000000", -- ADI R5,R7,0
	B"0101_000_110_000000",	--SW R0,R6,0
    others => X"FFFF") ;
begin

    data_out <= memory(to_integer(unsigned(address)));

end arc_Imem;

